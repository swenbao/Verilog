module top();

input clk, reset, in;
wire clock_div, tmp;
